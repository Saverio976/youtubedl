module youtubedl

pub struct DownloadInfo {
pub:
	title string
	download_url string
	extension string
	length_seconds int
}
