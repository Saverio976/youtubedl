module youtubedl
